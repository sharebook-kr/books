`timescale 1ns/10ps 

module testbench;

initial begin
    $display("hello world");
end

endmodule